// Copyright 2023 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51

// gives us the `FF(...) macro making it easy to have properly defined flip-flops
`include "common_cells/registers.svh"

// simple ROM
module bootrom #(
  /// The OBI configuration for all ports.
  parameter obi_pkg::obi_cfg_t           ObiCfg      = obi_pkg::ObiDefaultConfig,
  /// The request struct.
  parameter type                         obi_req_t   = logic,
  /// The response struct.
  parameter type                         obi_rsp_t   = logic,

  /// Boot ROM base address
  parameter int                          BaseAddr = 32'h0300_D000,
  /// Boot ROM size in bytes
  parameter int                          SizeBytes = 'h1000
) (
  /// Clock
  input  logic clk_i,
  /// Active-low reset
  input  logic rst_ni,

  /// OBI request interface
  input  obi_req_t obi_req_i,
  /// OBI response interface
  output obi_rsp_t obi_rsp_o
);
  localparam int AddressLSB = 2; // LSB offset (2 bits for the byte address)
  localparam int SizeWords = SizeBytes >> AddressLSB; // Size in words
  localparam int SizeWordsLog2 = $clog2(SizeWords); // Size in words log2
  localparam int AddressMSB = SizeWordsLog2 + AddressLSB; // Address MSB (2 bits for the byte address)

  // Define some registers to hold the requests fields
  logic req_d, req_q; // Request valid
  logic we_d, we_q; // Write enable
  logic [ObiCfg.AddrWidth-1:0] addr_d, addr_q; // Internal address of the word to read
  logic [ObiCfg.IdWidth-1:0] id_d, id_q; // Id of the request, must be same for the response

  // Signals used to create the response
  logic [ObiCfg.DataWidth-1:0] rsp_data; // Data field of the obi response
  logic rsp_err; // Error field of the obi response

  // Wire the registers holding the request
  assign req_d = obi_req_i.req;
  assign id_d = obi_req_i.a.aid;
  assign we_d = obi_req_i.a.we;
  assign addr_d = obi_req_i.a.addr;
  always_ff @(posedge (clk_i) or negedge (rst_ni)) begin
    if (!rst_ni) begin
      req_q <= '0;
      id_q <= '0;
      we_q <= '0;
      addr_q <= '0;
    end else begin
      req_q <= req_d;
      id_q <= id_d;
      we_q <= we_d;
      addr_q <= addr_d;
    end
  end

  logic [ObiCfg.AddrWidth-1:0] addr_q_offset = addr_q - BaseAddr;

  // Full-width checks:
  //   misaligned    = any low 2 bits non-zero
  //   out_of_range  = any high bits above MSB set (i.e. addr_q >= size in bytes (SizeWords*4))
  logic misaligned = |addr_q_offset[AddressLSB-1:0];
  logic out_of_bounds = |addr_q_offset[ObiCfg.AddrWidth-1:AddressMSB];

  // Assign the response data
  logic [SizeWordsLog2-1:0] word_addr = addr_q_offset[AddressMSB-1:AddressLSB];

  always_comb begin
    rsp_data = '0;
    rsp_err  = '0;

    if(req_q) begin
      if(we_q) begin
        // $display(">> Boot ROM: write access: addr_q_offset = 0x%0h", addr_q_offset);
        // rsp_err = '1;
      end else if (misaligned || out_of_bounds) begin
        // $display(">> Boot ROM: misaligned or out of bounds access: addr_q = 0x%0h", addr_q_offset);
        rsp_err = '1;
      end else begin
        // $display(">> Boot ROM: read access: addr_q_offset = 0x%0h", addr_q_offset);
        rsp_data = rom_data[word_addr];
      end
    end
  end

  // Wire the response
  // A channel
  assign obi_rsp_o.gnt = obi_req_i.req;
  // R channel:
  assign obi_rsp_o.rvalid = req_q;
  assign obi_rsp_o.r.rdata = rsp_data;
  assign obi_rsp_o.r.rid = id_q;
  assign obi_rsp_o.r.err = rsp_err;
  assign obi_rsp_o.r.r_optional = '0;

  // Static ROM data
  logic [31:0] rom_data [0:SizeWords-1] = {
    // --- ROM STATIC DATA START ---
    32'h0CFF3197, 32'h00018193, 32'h0CFF3117, 32'h7F810113, // 0x0000 - 0x0003
    32'h00000297, 32'h57E28293, 32'h00018313, 32'h00018393, // 0x0004 - 0x0007
    32'h00730C63, 32'h0002AE03, 32'h01C32023, 32'h00428293, // 0x0008 - 0x000B
    32'h00430313, 32'hFEDFF06F, 32'h00018293, 32'h00018313, // 0x000C - 0x000F
    32'h00628863, 32'h0002A023, 32'h00428293, 32'hFF5FF06F, // 0x0010 - 0x0013
    32'h00000093, 32'h00000213, 32'h00000293, 32'h00000313, // 0x0014 - 0x0017
    32'h00000393, 32'h00000413, 32'h00000493, 32'h00000513, // 0x0018 - 0x001B
    32'h00000593, 32'h00000613, 32'h00000693, 32'h00000713, // 0x001C - 0x001F
    32'h00000793, 32'h204000EF, 32'hFFFF3297, 32'hF8028293, // 0x0020 - 0x0023
    32'h00A2A023, 32'h10500073, 32'hFA010113, 32'h04F12A23, // 0x0024 - 0x0027
    32'h04410793, 32'h02912A23, 32'h03212823, 32'h03312623, // 0x0028 - 0x002B
    32'h03412423, 32'h03512223, 32'h02112E23, 32'h02812C23, // 0x002C - 0x002F
    32'h03612023, 32'h01712E23, 32'h00050493, 32'h04B12223, // 0x0030 - 0x0033
    32'h04C12423, 32'h04D12623, 32'h04E12823, 32'h05012C23, // 0x0034 - 0x0037
    32'h05112E23, 32'h00F12023, 32'h02500913, 32'h07800993, // 0x0038 - 0x003B
    32'h06300A13, 32'h07300A93, 32'h0004C503, 32'h02051863, // 0x003C - 0x003F
    32'h03C12083, 32'h03812403, 32'h03412483, 32'h03012903, // 0x0040 - 0x0043
    32'h02C12983, 32'h02812A03, 32'h02412A83, 32'h02012B03, // 0x0044 - 0x0047
    32'h01C12B83, 32'h06010113, 32'h00008067, 32'h0D251863, // 0x0048 - 0x004B
    32'h0014C783, 32'h09379263, 32'h00012783, 32'h03000513, // 0x004C - 0x004F
    32'h00478713, 32'h00E12023, 32'h0007A703, 32'h08070063, // 0x0050 - 0x0053
    32'h00000413, 32'h00900593, 32'h00410B13, 32'h00F77793, // 0x0054 - 0x0057
    32'h00078613, 32'h00F5B7B3, 32'h40F007B3, 32'h0077F793, // 0x0058 - 0x005B
    32'h03078793, 32'h00F60633, 32'h008B06B3, 32'h00C68023, // 0x005C - 0x005F
    32'h00475713, 32'h00140793, 32'h02071463, 32'hFFF00B93, // 0x0060 - 0x0063
    32'h008B07B3, 32'h0007C503, 32'hFFF40413, 32'h0E8000EF, // 0x0064 - 0x0067
    32'hFF7418E3, 32'h00148493, 32'h00148493, 32'hF4DFF06F, // 0x0068 - 0x006B
    32'h00078413, 32'hFA9FF06F, 32'h01479E63, 32'h00012783, // 0x006C - 0x006F
    32'h0007C503, 32'h00478713, 32'h00E12023, 32'h0B8000EF, // 0x0070 - 0x0073
    32'hFD5FF06F, 32'hFD5798E3, 32'h00012783, 32'h0007A403, // 0x0074 - 0x0077
    32'h00478713, 32'h00E12023, 32'h00044503, 32'hFA050CE3, // 0x0078 - 0x007B
    32'h00140413, 32'h090000EF, 32'hFF1FF06F, 32'h088000EF, // 0x007C - 0x007F
    32'hFA9FF06F, 32'h03002737, 32'h00070223, 32'hF8000693, // 0x0080 - 0x0083
    32'h00D70623, 32'h00A00613, 32'h00C70023, 32'h00070793, // 0x0084 - 0x0087
    32'h00070223, 32'h00300713, 32'h00E78623, 32'hFC700713, // 0x0088 - 0x008B
    32'h00E78423, 32'h02000713, 32'h00E78823, 32'h00008067, // 0x008C - 0x008F
    32'h03002737, 32'h01470713, 32'h00074783, 32'h0207F793, // 0x0090 - 0x0093
    32'hFE078CE3, 32'h030027B7, 32'h00A78023, 32'h00008067, // 0x0094 - 0x0097
    32'h030027B7, 32'h01478793, 32'h0007C703, 32'h02077713, // 0x0098 - 0x009B
    32'hFE070CE3, 32'h0007C703, 32'h04077713, 32'hFE0706E3, // 0x009C - 0x009F
    32'h00008067, 32'hFBDFF06F, 32'hFF010113, 32'h200107B7, // 0x00A0 - 0x00A3
    32'h00112623, 32'h00812423, 32'h00912223, 32'h0007A023, // 0x00A4 - 0x00A7
    32'hF65FF0EF, 32'h00000517, 32'h1DC50513, 32'hDEDFF0EF, // 0x00A8 - 0x00AB
    32'h10000437, 32'hFADFF0EF, 32'h10042783, 32'h00178793, // 0x00AC - 0x00AF
    32'h10F42023, 32'h10042703, 32'h00300793, 32'h00E7FE63, // 0x00B0 - 0x00B3
    32'h00000517, 32'h1C050513, 32'h10040413, 32'hDBDFF0EF, // 0x00B4 - 0x00B7
    32'hF81FF0EF, 32'h00042023, 32'h100007B7, 32'h1007A703, // 0x00B8 - 0x00BB
    32'h00300493, 32'h10078793, 32'h04971A63, 32'h00000517, // 0x00BC - 0x00BF
    32'h1B450513, 32'hD95FF0EF, 32'h03000437, 32'hF55FF0EF, // 0x00C0 - 0x00C3
    32'h01842583, 32'h00000517, 32'h1D050513, 32'hD7DFF0EF, // 0x00C4 - 0x00C7
    32'hF41FF0EF, 32'h01842783, 32'h00078293, 32'h00028067, // 0x00C8 - 0x00CB
    32'h00050593, 32'h00000517, 32'h1C850513, 32'hD5DFF0EF, // 0x00CC - 0x00CF
    32'hF21FF0EF, 32'h10500073, 32'hFFDFF06F, 32'h0007A583, // 0x00D0 - 0x00D3
    32'h00000517, 32'h1D050513, 32'h20010437, 32'h00158593, // 0x00D4 - 0x00D7
    32'hD39FF0EF, 32'hEFDFF0EF, 32'h600007B7, 32'hFE87A783, // 0x00D8 - 0x00DB
    32'h02000713, 32'h600007B7, 32'hFFC7A783, 32'h00000517, // 0x00DC - 0x00DF
    32'h1B450513, 32'h600007B7, 32'hFF87A783, 32'h600007B7, // 0x00E0 - 0x00E3
    32'hFF47A783, 32'h600007B7, 32'hFF07A783, 32'h600007B7, // 0x00E4 - 0x00E7
    32'hFEC7A783, 32'h600007B7, 32'hFEE7A023, 32'hCEDFF0EF, // 0x00E8 - 0x00EB
    32'hEB1FF0EF, 32'h600007B7, 32'h00942023, 32'h0007A783, // 0x00EC - 0x00EF
    32'h00000517, 32'h18850513, 32'h600007B7, 32'h2007A783, // 0x00F0 - 0x00F3
    32'h600007B7, 32'h4007A783, 32'h600007B7, 32'h6007A783, // 0x00F4 - 0x00F7
    32'h600017B7, 32'h8007A783, 32'h600017B7, 32'hA007A783, // 0x00F8 - 0x00FB
    32'h600017B7, 32'hC007A783, 32'h600017B7, 32'hE007A783, // 0x00FC - 0x00FF
    32'h600017B7, 32'h0007A783, 32'h600017B7, 32'h2007A783, // 0x0100 - 0x0103
    32'h600017B7, 32'h4007A783, 32'h600017B7, 32'h6007A783, // 0x0104 - 0x0107
    32'hC79FF0EF, 32'hE3DFF0EF, 32'h00100793, 32'h00F42023, // 0x0108 - 0x010B
    32'h00000517, 32'h12C50513, 32'hC61FF0EF, 32'h03000437, // 0x010C - 0x010F
    32'hE21FF0EF, 32'h01C42583, 32'h00000517, 32'h09C50513, // 0x0110 - 0x0113
    32'hC49FF0EF, 32'hE0DFF0EF, 32'h01C42783, 32'h00078293, // 0x0114 - 0x0117
    32'h00028067, 32'h00050593, 32'h00000517, 32'h10050513, // 0x0118 - 0x011B
    32'hC29FF0EF, 32'hDEDFF0EF, 32'h10500073, 32'hFFDFF06F, // 0x011C - 0x011F
    32'h3E3E5242, 32'h61745320, 32'h64657472, 32'h0000000A, // 0x0120 - 0x0123
    32'h3E3E5242, 32'h73655220, 32'h69747465, 32'h7220676E, // 0x0124 - 0x0127
    32'h79727465, 32'h756F6320, 32'h7265746E, 32'h0000000A, // 0x0128 - 0x012B
    32'h3E3E5242, 32'h6F6F5420, 32'h6E616D20, 32'h65722079, // 0x012C - 0x012F
    32'h65697274, 32'h73202C73, 32'h7070696B, 32'h20676E69, // 0x0130 - 0x0133
    32'h74696E69, 32'h696C6169, 32'h6974617A, 32'h0A216E6F, // 0x0134 - 0x0137
    32'h00000000, 32'h3E3E5242, 32'h6D754A20, 32'h676E6970, // 0x0138 - 0x013B
    32'h206F7420, 32'h78257830, 32'h0000000A, 32'h3E3E5242, // 0x013C - 0x013F
    32'h74655220, 32'h206E7275, 32'h756C6176, 32'h72662065, // 0x0140 - 0x0143
    32'h53206D6F, 32'h3A4D4152, 32'h25783020, 32'h00000A78, // 0x0144 - 0x0147
    32'h3E3E5242, 32'h79725420, 32'h0A782520, 32'h00000000, // 0x0148 - 0x014B
    32'h3E3E5242, 32'h50535420, 32'h6E692049, 32'h61697469, // 0x014C - 0x014F
    32'h657A696C, 32'h00000A64, 32'h3E3E5242, 32'h6F6C4220, // 0x0150 - 0x0153
    32'h20736B63, 32'h64616F6C, 32'h000A6465, 32'h3E3E5242, // 0x0154 - 0x0157
    32'h6E6F4420, 32'h000A2165, 32'h3E3E5242, 32'h74655220, // 0x0158 - 0x015B
    32'h206E7275, 32'h756C6176, 32'h72662065, 32'h53206D6F, // 0x015C - 0x015F
    32'h61432044, 32'h203A6472, 32'h78257830, 32'h0000000A, // 0x0160 - 0x0163
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0164 - 0x0167
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0168 - 0x016B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x016C - 0x016F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0170 - 0x0173
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0174 - 0x0177
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0178 - 0x017B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x017C - 0x017F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0180 - 0x0183
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0184 - 0x0187
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0188 - 0x018B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x018C - 0x018F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0190 - 0x0193
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0194 - 0x0197
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0198 - 0x019B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x019C - 0x019F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01A0 - 0x01A3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01A4 - 0x01A7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01A8 - 0x01AB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01AC - 0x01AF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01B0 - 0x01B3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01B4 - 0x01B7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01B8 - 0x01BB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01BC - 0x01BF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01C0 - 0x01C3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01C4 - 0x01C7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01C8 - 0x01CB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01CC - 0x01CF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01D0 - 0x01D3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01D4 - 0x01D7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01D8 - 0x01DB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01DC - 0x01DF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01E0 - 0x01E3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01E4 - 0x01E7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01E8 - 0x01EB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01EC - 0x01EF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01F0 - 0x01F3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01F4 - 0x01F7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01F8 - 0x01FB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x01FC - 0x01FF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0200 - 0x0203
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0204 - 0x0207
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0208 - 0x020B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x020C - 0x020F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0210 - 0x0213
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0214 - 0x0217
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0218 - 0x021B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x021C - 0x021F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0220 - 0x0223
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0224 - 0x0227
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0228 - 0x022B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x022C - 0x022F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0230 - 0x0233
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0234 - 0x0237
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0238 - 0x023B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x023C - 0x023F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0240 - 0x0243
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0244 - 0x0247
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0248 - 0x024B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x024C - 0x024F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0250 - 0x0253
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0254 - 0x0257
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0258 - 0x025B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x025C - 0x025F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0260 - 0x0263
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0264 - 0x0267
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0268 - 0x026B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x026C - 0x026F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0270 - 0x0273
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0274 - 0x0277
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0278 - 0x027B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x027C - 0x027F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0280 - 0x0283
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0284 - 0x0287
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0288 - 0x028B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x028C - 0x028F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0290 - 0x0293
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0294 - 0x0297
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0298 - 0x029B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x029C - 0x029F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02A0 - 0x02A3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02A4 - 0x02A7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02A8 - 0x02AB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02AC - 0x02AF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02B0 - 0x02B3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02B4 - 0x02B7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02B8 - 0x02BB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02BC - 0x02BF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02C0 - 0x02C3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02C4 - 0x02C7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02C8 - 0x02CB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02CC - 0x02CF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02D0 - 0x02D3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02D4 - 0x02D7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02D8 - 0x02DB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02DC - 0x02DF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02E0 - 0x02E3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02E4 - 0x02E7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02E8 - 0x02EB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02EC - 0x02EF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02F0 - 0x02F3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02F4 - 0x02F7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02F8 - 0x02FB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x02FC - 0x02FF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0300 - 0x0303
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0304 - 0x0307
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0308 - 0x030B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x030C - 0x030F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0310 - 0x0313
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0314 - 0x0317
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0318 - 0x031B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x031C - 0x031F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0320 - 0x0323
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0324 - 0x0327
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0328 - 0x032B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x032C - 0x032F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0330 - 0x0333
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0334 - 0x0337
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0338 - 0x033B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x033C - 0x033F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0340 - 0x0343
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0344 - 0x0347
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0348 - 0x034B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x034C - 0x034F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0350 - 0x0353
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0354 - 0x0357
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0358 - 0x035B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x035C - 0x035F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0360 - 0x0363
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0364 - 0x0367
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0368 - 0x036B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x036C - 0x036F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0370 - 0x0373
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0374 - 0x0377
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0378 - 0x037B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x037C - 0x037F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0380 - 0x0383
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0384 - 0x0387
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0388 - 0x038B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x038C - 0x038F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0390 - 0x0393
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0394 - 0x0397
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x0398 - 0x039B
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x039C - 0x039F
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03A0 - 0x03A3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03A4 - 0x03A7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03A8 - 0x03AB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03AC - 0x03AF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03B0 - 0x03B3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03B4 - 0x03B7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03B8 - 0x03BB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03BC - 0x03BF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03C0 - 0x03C3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03C4 - 0x03C7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03C8 - 0x03CB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03CC - 0x03CF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03D0 - 0x03D3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03D4 - 0x03D7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03D8 - 0x03DB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03DC - 0x03DF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03E0 - 0x03E3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03E4 - 0x03E7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03E8 - 0x03EB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03EC - 0x03EF
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03F0 - 0x03F3
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03F4 - 0x03F7
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, // 0x03F8 - 0x03FB
    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000 // 0x03FC - 0x03FF
    // --- ROM STATIC DATA END ---
  };

endmodule